package package_dpram;
	`include "transaction.sv"
	`include "packet_generator.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "scoreboard.sv"
	`include "environment.sv"
	`include "test.sv"
endpackage

