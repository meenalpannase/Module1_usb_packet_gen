//`ifdef defines.sv
//Calling the DUT

//Calling the DPRAM package

//Calling the interface

//Calling the test

//Calling the scoreboard

module top();
	//Importing the DPRAM package
	
 	//Declaring variables for clock and reset
 	
	//Generating the clock
 	
	//Instantiating the interface
 
	//Calling the DUT
	
		
	//Calling the test
	
	//Calling the run task to start the testbench execution	
	initial 
	begin
		
	end
endmodule
//`endif
