`ifdef defines.sv
//Include the transaction

class scoreboard;
	//Transaction class handle
	
	//Mailbox for driver to scoreboard
	
	//Mailbox from monitor to scoreboard
	
	//2-D Array for storing data from driver and monitor
	
	//Variables to indicates the status
	
	
	//Connecting driver and scoreboard, monitor and scoreboard with mailboc
	

	//Task to collect data from driver and monitor and store them in memories
	
				//Getting the driver transaction from mailbox		
				
			
				//Getting the monitor transaction from mailbox		
				
	endtask
	
	//Task to compare memories and generate report
	
endclass
`endif
