#`timescale 
#`define DATA_WIDTH 
#`define ADDR_WIDTH 
#`define DATA_DEPTH 
