`ifdef defines.sv
//Calling the transaction_DPRAM

class generator;
	//Transcation handle
	
	//Mailbox for generator to driver connection
	

	//Function to connect generator and driver using mailbox
	

	//Creating a task to generate the random stimuli
	
`endif
endclass
