`timescale 1ns/100ps
`define DATA_WIDTH 128
`define ADDR_WIDTH 16
`define DATA_DEPTH 65536
