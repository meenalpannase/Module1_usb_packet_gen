//`ifdef defines.sv
//Including the environment

class test;
	//Virtual interfaces for driver and monitor
 	
 	//environment handle
 	
 	
	//Function to connect the virtual interfaces from driver and monitor to test
 	
	//Task to start the methods of the environment
 	
endclass
//`endif
