package package_dpram;
	
endpackage

