//`ifdef defines.sv
//Calling the transaction class

class monitor;
	//Transaction handle

	//Mailbox from monitor to scoreboard
	
	//Virtual interfacewith monitor modport
	

	//Functional coverage for outputs
	

	//Function to connect the monitor and scoreboard with mailbox and virtual interface from driver to environmnet
	
	//Creating object for covergroup
		
	//Task to collect output from interface
	
endclass
`endif
