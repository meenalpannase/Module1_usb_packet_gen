`ifdef defines.sv
class transaction;
	//Randomizing input variables
	
	//Output variable declaration
	

	//Copying objects to run different test cases using same transaction class
	
endclass
`endif
