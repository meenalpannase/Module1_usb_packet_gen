`ifdef defines.sv
//Calling the packet generator

//Calling the transaction class

class driver
	//transaction class handle
	
	//Mailbox for generator to driver connection
	
	//Mailbox for driver to scoreboard connection

	//Virtual interface
	

	//Functional coverage for inputs
	

	//Function to connect the driver and generator, driver to scoreboard with mailbox and virtual interface 	//from driver to environmnet
	

	//Task to drive the stimulus
	
				//Put randomized inputs in mailbox from driver to scoreboard			
				
				//Covergroup sampling
				
				
			
	
endclass
`endif
